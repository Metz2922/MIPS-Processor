library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

  

entity barrelshifter is
port 	(data_in : in std_logic_vector(31 downto 0);
	 ctrl	: in std_logic_vector(4 downto 0);
	 typesel: in std_logic; --Logical when 0 arithmetic when 1
	 rlsel:   in std_logic; --Shifts right when 0 left when 1
	 data_out : out std_logic_vector(31 downto 0));
end barrelshifter;




architecture mixed of barrelshifter is





component mux2t1_N is
  generic(N : integer := 32); -- Generic of type integer for input/output data width. Default value is 32.
  port(i_S          : in std_logic;
       i_D0         : in std_logic_vector(N-1 downto 0);
       i_D1         : in std_logic_vector(N-1 downto 0);
       o_O          : out std_logic_vector(N-1 downto 0));

end component;

component mux2t1d is
  port(i_S          : in std_logic;
       i_D0         : in std_logic;
       i_D1         : in std_logic;
       o_O          : out std_logic);

end component;

signal mux4to3	: std_logic_vector(31 downto 0);
signal mux3to2	: std_logic_vector(31 downto 0);
signal mux2to1	: std_logic_vector(31 downto 0);
signal mux1to0	: std_logic_vector(31 downto 0);
signal D1	: std_logic;
signal D1_ext	: std_logic_vector(31 downto 0);
signal invdata : std_logic_vector(31 downto 0);
signal muxdatain : std_logic_vector(31 downto 0);
signal invdataout : std_logic_vector(31 downto 0);
signal data	: std_logic_vector(31 downto 0);
begin


gen: for i in 0 to 31 generate
invdata(31-i) <= data_in(i);
end generate;


muxAorL: mux2t1d port map(
	i_S => typesel,
	i_D0 => '0',
	i_D1 => data_in(31),
	o_O => D1);


muxRorLin: mux2t1_N port map(
	i_S => rlsel,
	i_D0 => data_in,
	i_D1 => invdata,
	o_O => muxdatain);

D1_ext <= (31 downto 0 => D1);




  l4ext: for i in 31 downto 16 generate
    MUXI: mux2t1d port map(
              i_S      => ctrl(4),      
              i_D0     => muxdatain(i),  
              i_D1     => D1,
              o_O      => mux4to3(i)); 
  end generate l4ext;
  
    l4data: for i in 15 downto 0 generate
    MUXI: mux2t1d port map(
              i_S      => ctrl(4),      
              i_D0     => muxdatain(i),  
              i_D1     => muxdatain(i+16),
              o_O      => mux4to3(i)); 
  end generate l4data;
  

   l3ext: for i in 31 downto 24 generate
    MUXI: mux2t1d port map(
              i_S      => ctrl(3),      
              i_D0     => mux4to3(i),  
              i_D1     => D1,
              o_O      => mux3to2(i)); 
  end generate l3ext;
  
    l3data: for i in 23 downto 0 generate
    MUXI: mux2t1d port map(
              i_S      => ctrl(3),      
              i_D0     => mux4to3(i),  
              i_D1     => mux4to3(i+8),
              o_O      => mux3to2(i)); 
  end generate l3data;
  
   l2ext: for i in 31 downto 28 generate
    MUXI: mux2t1d port map(
              i_S      => ctrl(2),      
              i_D0     => mux3to2(i),  
              i_D1     => D1,
              o_O      => mux2to1(i)); 
  end generate l2ext;
  
    l2data: for i in 27 downto 0 generate
    MUXI: mux2t1d port map(
              i_S      => ctrl(2),      
              i_D0     => mux3to2(i),  
              i_D1     => mux3to2(i+4),
              o_O      => mux2to1(i)); 
  end generate l2data;
  

   l1ext: for i in 31 downto 30 generate
    MUXI: mux2t1d port map(
              i_S      => ctrl(1),      
              i_D0     => mux2to1(i),  
              i_D1     => D1,
              o_O      => mux1to0(i)); 
  end generate l1ext;
  
    l1data: for i in 29 downto 0 generate
    MUXI: mux2t1d port map(
              i_S      => ctrl(1),      
              i_D0     => mux2to1(i),  
              i_D1     => mux2to1(i+2),
              o_O      => mux1to0(i)); 
  end generate l1data;





    l0ext: mux2t1d port map(
              i_S      => ctrl(0),      
              i_D0     => mux1to0(31),  
              i_D1     => D1,
              o_O      => data(31)); 

  
    l0data: for i in 30 downto 0 generate
    MUXI: mux2t1d port map(
              i_S      => ctrl(0),      
              i_D0     => mux1to0(i),  
              i_D1     => mux1to0(i+1),
              o_O      => data(i)); 
  end generate l0data;


gen2: for i in 0 to 31 generate
invdataout(31-i) <= data(i);
end generate;

muxRorLout: mux2t1_N port map(
	i_S => rlsel,
	i_D0 => data,
	i_D1 => invdataout,
	o_O => data_out);





end mixed;