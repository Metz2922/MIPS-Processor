library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ALU is
port(	i_A	: in std_logic_vector(31 downto 0);
	i_B	: in std_logic_vector(31 downto 0);
	i_ALUc	: in std_logic_vector(6 downto 0);
	i_shamt	: in std_logic_vector(4 downto 0);
	i_signed: in std_logic;
	i_replimm : in std_logic_vector(7 downto 0);
	o_Zero	: out std_logic;
	o_O	: out std_logic_vector(31 downto 0);
	o_C	: out std_logic;
	o_Ovf	: out std_logic);
end ALU;
	



architecture structural of ALU is

component nAdd_Sub is
	generic(N : integer := 32);
	port(i_A	: in std_logic_vector(N-1 downto 0);
		i_B	: in std_logic_vector(N-1 downto 0);
		i_CTRL	: in std_logic;
		o_S	: out std_logic_vector(N-1 downto 0);
		o_C	: out std_logic;
		o_Ovf	: out std_logic);
end component;

component SLT is
port(i_D: in std_logic;
	o_D: out std_logic_vector(31 downto 0));
end component;

component barrelshifter is
port 	(data_in : in std_logic_vector(31 downto 0);
	 ctrl	: in std_logic_vector(4 downto 0);
	 typesel: in std_logic; --Logical when 0 arithmetic when 1
	 rlsel:   in std_logic; --Shifts right when 0 left when 1
	 data_out : out std_logic_vector(31 downto 0));
end component;

component zeroDetect is
port(i_D	: in std_logic_vector(31 downto 0);
	o_Z	: out std_logic);
end component;

component mux2t1_N is
  generic(N : integer := 16);
  port(i_S          : in std_logic;
       i_D0         : in std_logic_vector(N-1 downto 0);
       i_D1         : in std_logic_vector(N-1 downto 0);
       o_O          : out std_logic_vector(N-1 downto 0));
end component;

component onesComp is
	generic(N : integer := 32);
	port(i_D0	: in std_logic_vector(N-1 downto 0);
	o_F		: out std_logic_vector(N-1 downto 0));
end component;

component andgN is
	generic(N : integer := 32);
	port(i_D0	: in std_logic_vector(N-1 downto 0);
	i_D1		: in std_logic_vector(N-1 downto 0);
	o_F		: out std_logic_vector(N-1 downto 0));
end component;

component orgN is
	generic(N : integer := 32);
	port(i_D0	: in std_logic_vector(N-1 downto 0);
	i_D1		: in std_logic_vector(N-1 downto 0);
	o_F		: out std_logic_vector(N-1 downto 0));
end component;

component xorgN is
	generic(N : integer := 32);
	port(i_D0	: in std_logic_vector(N-1 downto 0);
	i_D1		: in std_logic_vector(N-1 downto 0);
	o_F		: out std_logic_vector(N-1 downto 0));
end component;

signal s_O : std_logic_vector(31 downto 0);
signal s_AND, s_ADD, s_OR, s_NOR, s_XOR, s_BARR, s_SLT : std_logic_vector(31 downto 0);
signal s_BARRELCTRL : std_logic_vector(4 downto 0);
signal s_MUX5O : std_logic_vector(31 downto 0);
signal s_MUX4O, s_MUX3O, replout : std_logic_vector(31 downto 0);
signal s_MUX2O, s_MUX1O, s_mux0O : std_logic_vector(31 downto 0);
signal Overflow		: std_logic;

begin

replout <= i_replimm & i_replimm & i_replimm & i_replimm;

ANDG: andgN
port MAP(i_D0 =>  i_A,
	i_D1 => i_B,
	o_F => s_AND);

ADDER: nAdd_Sub
port MAP(i_A => i_B,-- its backwards
	i_B => i_A,
	i_CTRL => i_ALUc(3),
	o_S => s_ADD,
	o_C => o_C,
	o_Ovf => Overflow);

ZERO: zeroDetect
port MAP(i_D => s_O,
	o_Z => o_Zero);

ORG: orgN
port MAP(i_D0 => i_A,
	i_D1 => i_B,
	o_F => s_OR);

NORG: onesComp
port MAP(i_D0 => s_OR,
	o_F => s_NOR);

XORG: xorgN
port MAP(i_D0 => i_A,
	i_D1 => i_B,
	o_F => s_XOR);

BARRELCTRL: mux2t1_N
generic MAP(N => 5)
port MAP(i_D0 => i_shamt,
	i_D1 => "10000",
	i_S => i_ALUc(4),
	o_O => s_BARRELCTRL);

BARREL: barrelshifter
port MAP(data_in => i_B,
	 ctrl	=> s_BARRELCTRL,
	 typesel => i_ALUc(1),
	 rlsel => i_ALUc(0),
	 data_out => s_BARR);

SLTFILL: SLT
port MAP(i_D => s_ADD(31),
	o_D => s_SLT);

MUX5: mux2t1_N
generic MAP(N => 32)
port MAP(i_D0 => s_OR,
	i_D1 => s_NOR,
	i_S => i_ALUc(3),
	o_O => s_MUX5O);

MUX4: mux2t1_N
generic MAP(N => 32)
port MAP(i_D0 => s_MUX5O,
	i_D1 => s_XOR,
	i_S => i_ALUc(1),
	o_O => s_MUX4O);

MUX3: mux2t1_N
generic MAP(N => 32)
port MAP(i_D0 => s_AND,
	i_D1 => s_ADD,
	i_S => i_ALUc(1),
	o_O => s_MUX3O);

MUX2: mux2t1_N
generic MAP(N => 32)
port MAP(i_D0 => s_BARR,
	i_D1 => s_SLT,
	i_S => i_ALUc(3),
	o_O => s_MUX2O);

MUX1: mux2t1_N
generic MAP(N => 32)
port MAP(i_D0 => s_MUX3O,
	i_D1 => s_MUX4O,
	i_S => i_ALUc(0),
	o_O => s_MUX1O);

MUX0: mux2t1_N
generic MAP(N => 32)
port MAP(i_D0 => s_MUX1O,
	i_D1 => s_MUX2O,
	i_S => i_ALUc(2),
	o_O => s_MUX0O);

replMux: mux2t1_N
generic MAP(N => 32)
port MAP(i_D0 => s_MUX0O,
	i_D1 => replout,
	i_S => i_ALUc(6),
	o_O => s_O);


o_O <= s_O;
o_Ovf <= Overflow AND i_ALUc(5);
end structural;
