library IEEE;
use IEEE.std_logic_1164.all;
use work.bus_mux_input.all;
use IEEE.numeric_std.all;

entity tb_registerFile is
end tb_registerFile;

architecture mixed of tb_registerFile is

component registerFile is
	port(i_D: in std_logic_vector(31 downto 0);
		i_CLK: in std_logic;
		i_RST: in std_logic;
		i_DS: in std_logic_vector(4 downto 0);
		i_RS: in std_logic_vector(4 downto 0);
		i_RT: in std_logic_vector(4 downto 0);
		o_RS: out std_logic_vector(31 downto 0);
		o_RT: out std_logic_vector(31 downto 0);
		i_WE: in std_logic);
end component;

signal s_D, s_oRS, s_oRT: std_logic_vector(31 downto 0);
signal s_CLK, s_RST, s_WE: std_logic;
signal s_DS, s_iRS, s_iRT: std_logic_vector(4 downto 0);

begin

DUT0: registerFile
port MAP(i_D => s_D,
	i_CLK => s_CLK,
	i_RST => s_RST,
	i_DS => s_DS,
	i_RS => s_iRS,
	i_RT => s_iRT,
	o_RS => s_oRS,
	o_RT => s_oRT,
	i_WE => s_WE);

P_CLK: process
begin
	s_CLK <= '1';
	wait for 10 ns;
	s_CLK <= '0';
	wait for 10 ns;
end process;

P_TESTS: process
begin
	s_RST <= '1';
	wait for 10 ns;
	s_RST <= '0';
	wait for 10 ns;

	s_iRS <= "00000";
	s_iRT <= "00000";
	wait for 10 ns;
	
	s_DS <= "00001";
	s_D <= "11111111111111111111111111111111";
	s_iRS <= "00001";
	s_WE <= '1';
	wait for 10 ns;

	s_DS <= "00000";
	s_WE <= '0';
	wait for 10 ns;

	s_DS <= "00111";
	s_D <= "10101011010110101011010110101011";
	s_WE <= '1';
	wait for 10 ns;
	
	s_DS <= "00000";
	s_iRT <= "00111";
	s_WE <= '0';
	wait for 10 ns;

	wait for 10 ns;

end process;
end mixed;
