library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tb_PC is
end tb_PC;

architecture mixed of tb_PC is

component PC is
port(i_CLK	: in std_logic;
	i_RST	: in std_logic;
	i_CHANGE: in std_logic_vector(31 downto 0); -- Drop in program counter
	o_PC	: out std_logic_vector(31 downto 0)); -- To read input of instruction mem
end component;

signal s_CLK, s_RST : std_logic;
signal s_CHANGE: std_logic_vector(31 downto 0);
signal s_PC: std_logic_vector(31 downto 0);

begin

DUT0: PC
port MAP(i_CLK => s_CLK,
	i_CHANGE => s_CHANGE,
	i_RST => s_RST,
	o_PC => s_PC);

P_CLK: process
begin
	s_CLK <= '1';
	wait for 10 ns;
	s_CLK <= '0';
	wait for 10 ns;
end process;

P_TESTS: process
begin
	s_RST <= '0';
	s_CHANGE <= x"00000000";
	wait for 50 ns;

	s_CHANGE <= x"00010C00";
	wait for 20 ns;

	s_CHANGE <= x"00A1011C";
	wait for 40 ns;
	
	s_CHANGE <= x"00A10120";
	wait for 10 ns;

	s_CHANGE <= x"00A10124";
	wait for 10 ns;

	s_RST <= '1';
	wait for 10 ns;

end process;
end mixed;
