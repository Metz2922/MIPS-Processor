library IEEE;
use IEEE.std_logic_1164.all;

entity nAdd_Sub is
	generic(N : integer := 32);
	port(i_A	: in std_logic_vector(N-1 downto 0);
		i_B	: in std_logic_vector(N-1 downto 0);
		i_CTRL	: in std_logic;
		o_S	: out std_logic_vector(N-1 downto 0);
		o_C	: out std_logic;
		o_Ovf	: out std_logic);
end nAdd_Sub;

architecture structural of nAdd_Sub is

component rippleAdder_N is
	generic(N : integer := 32);
	port(i_C	: in std_logic;
		i_A	: in std_logic_vector(N-1 downto 0);
		i_B	: in std_logic_vector(N-1 downto 0);
		o_O	: out std_logic_vector(N-1 downto 0);
		o_C	: out std_logic);
end component;

component onesComp is
	generic(N : integer := 32);
	port(i_D0	: in std_logic_vector(N-1 downto 0);
	o_F		: out std_logic_vector(N-1 downto 0));
end component;

component mux2t1_N is
generic(N : integer := 16);
port (i_S          : in std_logic;
       i_D0         : in std_logic_vector(N-1 downto 0);
       i_D1         : in std_logic_vector(N-1 downto 0);
       o_O          : out std_logic_vector(N-1 downto 0));
end component;

signal s_IA : std_logic_vector(N-1 downto 0);
signal s_muxA : std_logic_vector(N-1 downto 0);
signal s_OS : std_logic_vector(N-1 downto 0);

begin

invertA: onesComp
port MAP(i_D0 => i_A,
	o_F => s_IA);

muxA: mux2t1_N
generic MAP(N => 32)
port MAP(i_S => i_CTRL,
	i_D0 => i_A,
	i_D1 => s_IA,
	o_O => s_muxA);

adder: rippleAdder_N
port MAP(i_C => i_CTRL,
	i_A => s_muxA,
	i_B => i_B,
	o_O => s_OS,
	o_C => o_C);

--o_Ovf <= o_C AND i_CTRL;
o_Ovf <= (NOT s_muxA(N-1) AND NOT i_B(N-1) AND s_OS(N-1)) OR (s_muxA(N-1) AND i_B(N-1) AND NOT s_OS(N-1));
o_S <= s_OS;

end structural;
