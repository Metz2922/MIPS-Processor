library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity PC is
	port(i_CLK	: in std_logic;
		i_RST	: in std_logic;
		i_CHANGE: in std_logic_vector(31 downto 0); -- Drop in program counter
		WE		: in std_logic;
		o_PC	: out std_logic_vector(31 downto 0)); -- To read input of instruction mem
end PC;

architecture rtl of PC is
signal s_NEWVAL : std_logic_vector(31 downto 0);


begin
process(i_CLK)
begin
if(rising_edge(i_CLK)) then
	if(i_RST = '1') then
		s_NEWVAL <= x"00400000";
	else
		s_NEWVAL <= i_CHANGE;
	end if;
end if;
o_PC <= s_NEWVAL when WE else o_PC;
end process;

end rtl;
