library IEEE;
use IEEE.std_logic_1164.all;

entity orgN is
	generic(N : integer := 32);
	port(i_D0	: in std_logic_vector(N-1 downto 0);
	i_D1		: in std_logic_vector(N-1 downto 0);
	o_F		: out std_logic_vector(N-1 downto 0));

end orgN;

architecture structural of orgN is

component org2 is
	port(i_A          : in std_logic;
	i_B		: in std_logic;
	o_F          : out std_logic);
end component;

begin

G_NBit_ORG: for i in 0 to N-1 generate
ORI: org2 port map(
	i_A => i_D0(i),
	i_B => i_D1(i),
	o_F => o_F(i));
end generate G_NBit_ORG;

end structural;